library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_unsigned.all;

package const_def is 
        constant DATA_SIZE : integer :=64;
        constant KEY_SIZE  : integer :=128;
	constant WORD_SIZE : integer := 32;        
	constant WORDS_NB  : integer :=  4; 
	constant CONST_SEQU: integer :=  3;    
	constant NB_ROUND  : integer := 44;
end const_def;
